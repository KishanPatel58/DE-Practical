<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0,0,139.4,-83.8</PageViewport></page 0>
<page 1>
<PageViewport>0,0,139.4,-83.8</PageViewport></page 1>
<page 2>
<PageViewport>0,0,139.4,-83.8</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-83.8</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-83.8</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-83.8</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-83.8</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-83.8</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-83.8</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-83.8</PageViewport></page 9></circuit>
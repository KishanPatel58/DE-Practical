<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>87.8189,-160.266,166.066,-207.304</PageViewport>
<gate>
<ID>2</ID>
<type>AE_DFF_LOW</type>
<position>121.5,-38.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>2 </output>
<input>
<ID>clock</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3</ID>
<type>AE_DFF_LOW</type>
<position>130.5,-38.5</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>3 </output>
<input>
<ID>clock</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4</ID>
<type>AE_DFF_LOW</type>
<position>139,-38.5</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>4 </output>
<input>
<ID>clock</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5</ID>
<type>AE_DFF_LOW</type>
<position>147,-38.5</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>5 </output>
<input>
<ID>clock</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>116.5,-36.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>9</ID>
<type>GA_LED</type>
<position>126,-35</position>
<input>
<ID>N_in2</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>GA_LED</type>
<position>135,-35</position>
<input>
<ID>N_in2</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>GA_LED</type>
<position>143,-35</position>
<input>
<ID>N_in2</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>GA_LED</type>
<position>151,-36.5</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>BB_CLOCK</type>
<position>112.5,-39.5</position>
<output>
<ID>CLK</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>130.5,-31</position>
<gparam>LABEL_TEXT Shift Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>130.5,-46.5</position>
<gparam>LABEL_TEXT 3-bit Up Asynchronous Counter using T-FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>112,-50.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>29</ID>
<type>BB_CLOCK</type>
<position>110,-58</position>
<output>
<ID>CLK</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>33</ID>
<type>BE_JKFF_LOW_NT</type>
<position>119.5,-54.5</position>
<input>
<ID>J</ID>17 </input>
<input>
<ID>K</ID>17 </input>
<output>
<ID>Q</ID>18 </output>
<input>
<ID>clock</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>34</ID>
<type>BE_JKFF_LOW_NT</type>
<position>130.5,-54.5</position>
<input>
<ID>J</ID>17 </input>
<input>
<ID>K</ID>17 </input>
<output>
<ID>Q</ID>19 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>35</ID>
<type>BE_JKFF_LOW_NT</type>
<position>140.5,-54.5</position>
<input>
<ID>J</ID>17 </input>
<input>
<ID>K</ID>17 </input>
<output>
<ID>Q</ID>24 </output>
<input>
<ID>clock</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>43</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>117,-77</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>28 </input>
<input>
<ID>IN_2</ID>27 </input>
<input>
<ID>IN_3</ID>25 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>45</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>138.5,-77.5</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>37 </input>
<input>
<ID>IN_2</ID>36 </input>
<input>
<ID>IN_3</ID>35 </input>
<input>
<ID>IN_4</ID>34 </input>
<input>
<ID>IN_5</ID>32 </input>
<input>
<ID>IN_6</ID>30 </input>
<input>
<ID>IN_7</ID>29 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_TOGGLE</type>
<position>110.5,-73.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_TOGGLE</type>
<position>110.5,-79.5</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_TOGGLE</type>
<position>110.5,-75.5</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_TOGGLE</type>
<position>110.5,-77.5</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_TOGGLE</type>
<position>125.5,-72.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>125.5,-74.5</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_TOGGLE</type>
<position>125.5,-76.5</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>59</ID>
<type>AA_TOGGLE</type>
<position>125.5,-78.5</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_TOGGLE</type>
<position>125.5,-80.5</position>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_TOGGLE</type>
<position>125.5,-82.5</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_TOGGLE</type>
<position>125.5,-84.5</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>63</ID>
<type>AA_TOGGLE</type>
<position>125.5,-86.5</position>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>65</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>153,-55</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>19 </input>
<input>
<ID>IN_2</ID>18 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>131,-91</position>
<gparam>LABEL_TEXT 3-bit Down Asynchronous Counter using T-FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>BE_JKFF_LOW_NT</type>
<position>120,-99</position>
<input>
<ID>J</ID>40 </input>
<input>
<ID>K</ID>40 </input>
<output>
<ID>Q</ID>51 </output>
<input>
<ID>clock</ID>54 </input>
<output>
<ID>nQ</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>70</ID>
<type>BE_JKFF_LOW_NT</type>
<position>131,-99</position>
<input>
<ID>J</ID>40 </input>
<input>
<ID>K</ID>40 </input>
<output>
<ID>Q</ID>52 </output>
<input>
<ID>clock</ID>48 </input>
<output>
<ID>nQ</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>71</ID>
<type>BE_JKFF_LOW_NT</type>
<position>141,-99</position>
<input>
<ID>J</ID>40 </input>
<input>
<ID>K</ID>40 </input>
<output>
<ID>Q</ID>50 </output>
<input>
<ID>clock</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>75</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>153.5,-99.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>52 </input>
<input>
<ID>IN_2</ID>51 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 7</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>77</ID>
<type>DA_FROM</type>
<position>112.5,-99</position>
<input>
<ID>IN_0</ID>54 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>81</ID>
<type>DE_TO</type>
<position>102.5,-99</position>
<input>
<ID>IN_0</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>83</ID>
<type>BB_CLOCK</type>
<position>95.5,-99</position>
<output>
<ID>CLK</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>85</ID>
<type>DE_TO</type>
<position>103.5,-95</position>
<input>
<ID>IN_0</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T</lparam></gate>
<gate>
<ID>87</ID>
<type>DA_FROM</type>
<position>108,-95</position>
<input>
<ID>IN_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T</lparam></gate>
<gate>
<ID>89</ID>
<type>AA_TOGGLE</type>
<position>99.5,-95</position>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>131.5,-112</position>
<gparam>LABEL_TEXT Mod-6 Asynchronous Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>BE_JKFF_LOW_NT</type>
<position>120.5,-120</position>
<input>
<ID>J</ID>70 </input>
<input>
<ID>K</ID>70 </input>
<output>
<ID>Q</ID>66 </output>
<input>
<ID>clear</ID>69 </input>
<input>
<ID>clock</ID>63 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>92</ID>
<type>BE_JKFF_LOW_NT</type>
<position>131.5,-120</position>
<input>
<ID>J</ID>71 </input>
<input>
<ID>K</ID>71 </input>
<output>
<ID>Q</ID>67 </output>
<input>
<ID>clear</ID>69 </input>
<input>
<ID>clock</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>93</ID>
<type>BE_JKFF_LOW_NT</type>
<position>141.5,-120</position>
<input>
<ID>J</ID>72 </input>
<input>
<ID>K</ID>72 </input>
<output>
<ID>Q</ID>68 </output>
<input>
<ID>clear</ID>69 </input>
<input>
<ID>clock</ID>67 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>95</ID>
<type>DA_FROM</type>
<position>113,-120</position>
<input>
<ID>IN_0</ID>63 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>96</ID>
<type>DE_TO</type>
<position>105,-120</position>
<input>
<ID>IN_0</ID>64 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>97</ID>
<type>BB_CLOCK</type>
<position>98,-120</position>
<output>
<ID>CLK</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>102</ID>
<type>BA_NAND2</type>
<position>153,-125</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>103</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>160,-130</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>67 </input>
<input>
<ID>IN_2</ID>66 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>105</ID>
<type>AA_TOGGLE</type>
<position>110.5,-116.5</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_TOGGLE</type>
<position>125,-116</position>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>107</ID>
<type>AA_TOGGLE</type>
<position>136,-116</position>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>108</ID>
<type>BE_JKFF_LOW_NT</type>
<position>120,-149.5</position>
<input>
<ID>J</ID>82 </input>
<input>
<ID>K</ID>82 </input>
<output>
<ID>Q</ID>86 </output>
<input>
<ID>clear</ID>78 </input>
<input>
<ID>clock</ID>73 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>109</ID>
<type>BE_JKFF_LOW_NT</type>
<position>131,-149.5</position>
<input>
<ID>J</ID>82 </input>
<input>
<ID>K</ID>82 </input>
<output>
<ID>Q</ID>87 </output>
<input>
<ID>clear</ID>78 </input>
<input>
<ID>clock</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>110</ID>
<type>BE_JKFF_LOW_NT</type>
<position>141,-149.5</position>
<input>
<ID>J</ID>82 </input>
<input>
<ID>K</ID>82 </input>
<output>
<ID>Q</ID>88 </output>
<input>
<ID>clear</ID>78 </input>
<input>
<ID>clock</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>111</ID>
<type>DA_FROM</type>
<position>112.5,-149.5</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cl</lparam></gate>
<gate>
<ID>112</ID>
<type>DE_TO</type>
<position>104.5,-149.5</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cl</lparam></gate>
<gate>
<ID>113</ID>
<type>BB_CLOCK</type>
<position>97.5,-149.5</position>
<output>
<ID>CLK</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>114</ID>
<type>BA_NAND2</type>
<position>152.5,-154.5</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>88 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>164.5,-159</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>90 </input>
<input>
<ID>IN_2</ID>91 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_TOGGLE</type>
<position>97.5,-143.5</position>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>119</ID>
<type>DE_TO</type>
<position>101.5,-143.5</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID TF</lparam></gate>
<gate>
<ID>120</ID>
<type>DA_FROM</type>
<position>109,-143</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID TF</lparam></gate>
<gate>
<ID>121</ID>
<type>DA_FROM</type>
<position>137,-138.5</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID QA</lparam></gate>
<gate>
<ID>122</ID>
<type>DE_TO</type>
<position>129.5,-138.5</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID QA</lparam></gate>
<gate>
<ID>123</ID>
<type>DA_FROM</type>
<position>146.5,-168</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID QB</lparam></gate>
<gate>
<ID>124</ID>
<type>DE_TO</type>
<position>139,-168</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID QB</lparam></gate>
<gate>
<ID>125</ID>
<type>DA_FROM</type>
<position>154.5,-164.5</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID QC</lparam></gate>
<gate>
<ID>126</ID>
<type>DE_TO</type>
<position>147,-164.5</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID QC</lparam></gate>
<gate>
<ID>128</ID>
<type>GA_LED</type>
<position>140,-138.5</position>
<input>
<ID>N_in0</ID>89 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>GA_LED</type>
<position>149.5,-168</position>
<input>
<ID>N_in0</ID>90 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>GA_LED</type>
<position>157.5,-164.5</position>
<input>
<ID>N_in0</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>133</ID>
<type>AA_LABEL</type>
<position>127,-173</position>
<gparam>LABEL_TEXT 3-bit Up Synchronous Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>BE_JKFF_LOW_NT</type>
<position>118.5,-188.5</position>
<input>
<ID>J</ID>97 </input>
<input>
<ID>K</ID>97 </input>
<output>
<ID>Q</ID>96 </output>
<input>
<ID>clock</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>136</ID>
<type>BE_JKFF_LOW_NT</type>
<position>130.5,-188.5</position>
<input>
<ID>J</ID>96 </input>
<input>
<ID>K</ID>96 </input>
<output>
<ID>Q</ID>94 </output>
<input>
<ID>clock</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>137</ID>
<type>BE_JKFF_LOW_NT</type>
<position>146,-189</position>
<input>
<ID>J</ID>95 </input>
<input>
<ID>K</ID>95 </input>
<output>
<ID>Q</ID>99 </output>
<input>
<ID>clock</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>141</ID>
<type>DE_TO</type>
<position>98.5,-188.5</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>143</ID>
<type>DA_FROM</type>
<position>111,-188.5</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>145</ID>
<type>BB_CLOCK</type>
<position>92.5,-188.5</position>
<output>
<ID>CLK</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>147</ID>
<type>AA_AND2</type>
<position>137,-181.5</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>149</ID>
<type>DE_TO</type>
<position>94,-184</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Switch</lparam></gate>
<gate>
<ID>151</ID>
<type>DA_FROM</type>
<position>110,-185</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Switch</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_TOGGLE</type>
<position>90,-184</position>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>155</ID>
<type>DE_TO</type>
<position>125.5,-183.5</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID qa</lparam></gate>
<gate>
<ID>156</ID>
<type>DE_TO</type>
<position>137,-185.5</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID qb</lparam></gate>
<gate>
<ID>157</ID>
<type>DE_TO</type>
<position>151.5,-182.5</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID qc</lparam></gate>
<gate>
<ID>158</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>160.5,-190</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>101 </input>
<input>
<ID>IN_2</ID>100 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 5</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>160</ID>
<type>DA_FROM</type>
<position>155.5,-189</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID qc</lparam></gate>
<gate>
<ID>162</ID>
<type>DA_FROM</type>
<position>154.5,-191.5</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID qb</lparam></gate>
<gate>
<ID>164</ID>
<type>DA_FROM</type>
<position>154.5,-194.5</position>
<input>
<ID>IN_0</ID>102 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID qa</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-36.5,118.5,-36.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-36.5,126,-36</points>
<connection>
<GID>9</GID>
<name>N_in2</name></connection>
<intersection>-36.5 1</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124.5,-36.5,127.5,-36.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-36.5,135,-36</points>
<connection>
<GID>11</GID>
<name>N_in2</name></connection>
<intersection>-36.5 1</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133.5,-36.5,136,-36.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-36.5,143,-36</points>
<connection>
<GID>12</GID>
<name>N_in2</name></connection>
<intersection>-36.5 1</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142,-36.5,144,-36.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>143 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-36.5,150,-36.5</points>
<connection>
<GID>13</GID>
<name>N_in0</name></connection>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-43.5,117.5,-39.5</points>
<intersection>-43.5 1</intersection>
<intersection>-39.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-43.5,144,-43.5</points>
<intersection>117.5 0</intersection>
<intersection>127.5 4</intersection>
<intersection>136 7</intersection>
<intersection>144 9</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116.5,-39.5,118.5,-39.5</points>
<connection>
<GID>2</GID>
<name>clock</name></connection>
<connection>
<GID>15</GID>
<name>CLK</name></connection>
<intersection>117.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>127.5,-43.5,127.5,-39.5</points>
<connection>
<GID>3</GID>
<name>clock</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>136,-43.5,136,-39.5</points>
<connection>
<GID>4</GID>
<name>clock</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>144,-43.5,144,-39.5</points>
<connection>
<GID>5</GID>
<name>clock</name></connection>
<intersection>-43.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-56.5,115,-49.5</points>
<intersection>-56.5 7</intersection>
<intersection>-52.5 8</intersection>
<intersection>-50.5 1</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114,-50.5,115,-50.5</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-49.5,135.5,-49.5</points>
<intersection>115 0</intersection>
<intersection>124.5 6</intersection>
<intersection>135.5 13</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>124.5,-56.5,124.5,-49.5</points>
<intersection>-56.5 10</intersection>
<intersection>-52.5 15</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>115,-56.5,116.5,-56.5</points>
<connection>
<GID>33</GID>
<name>K</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>115,-52.5,116.5,-52.5</points>
<connection>
<GID>33</GID>
<name>J</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>124.5,-56.5,127.5,-56.5</points>
<connection>
<GID>34</GID>
<name>K</name></connection>
<intersection>124.5 6</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>135.5,-56.5,135.5,-49.5</points>
<intersection>-56.5 17</intersection>
<intersection>-52.5 18</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>124.5,-52.5,127.5,-52.5</points>
<connection>
<GID>34</GID>
<name>J</name></connection>
<intersection>124.5 6</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>135.5,-56.5,137.5,-56.5</points>
<connection>
<GID>35</GID>
<name>K</name></connection>
<intersection>135.5 13</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>135.5,-52.5,137.5,-52.5</points>
<connection>
<GID>35</GID>
<name>J</name></connection>
<intersection>135.5 13</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>122.5,-63.5,148.5,-63.5</points>
<intersection>122.5 3</intersection>
<intersection>127.5 7</intersection>
<intersection>148.5 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>122.5,-63.5,122.5,-52.5</points>
<connection>
<GID>33</GID>
<name>Q</name></connection>
<intersection>-63.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>148.5,-63.5,148.5,-54</points>
<intersection>-63.5 1</intersection>
<intersection>-54 13</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>127.5,-63.5,127.5,-54.5</points>
<connection>
<GID>34</GID>
<name>clock</name></connection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>148.5,-54,150,-54</points>
<connection>
<GID>65</GID>
<name>IN_2</name></connection>
<intersection>148.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>134,-58.5,149,-58.5</points>
<intersection>134 3</intersection>
<intersection>136.5 8</intersection>
<intersection>149 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>134,-58.5,134,-52.5</points>
<intersection>-58.5 1</intersection>
<intersection>-52.5 9</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>149,-58.5,149,-55</points>
<intersection>-58.5 1</intersection>
<intersection>-55 11</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>136.5,-58.5,136.5,-54.5</points>
<intersection>-58.5 1</intersection>
<intersection>-54.5 10</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>133.5,-52.5,134,-52.5</points>
<connection>
<GID>34</GID>
<name>Q</name></connection>
<intersection>134 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>136.5,-54.5,137.5,-54.5</points>
<connection>
<GID>35</GID>
<name>clock</name></connection>
<intersection>136.5 8</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>149,-55,150,-55</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<intersection>149 7</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-58,114,-54.5</points>
<connection>
<GID>29</GID>
<name>CLK</name></connection>
<intersection>-54.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114,-54.5,116.5,-54.5</points>
<connection>
<GID>33</GID>
<name>clock</name></connection>
<intersection>114 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,-62.5,144.5,-52.5</points>
<intersection>-62.5 1</intersection>
<intersection>-52.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144.5,-62.5,150,-62.5</points>
<intersection>144.5 0</intersection>
<intersection>150 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>150,-62.5,150,-56</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>143.5,-52.5,144.5,-52.5</points>
<connection>
<GID>35</GID>
<name>Q</name></connection>
<intersection>144.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-75,114,-73.5</points>
<connection>
<GID>43</GID>
<name>IN_3</name></connection>
<intersection>-73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112.5,-73.5,114,-73.5</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>114 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-79.5,114,-78</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>-79.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112.5,-79.5,114,-79.5</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>114 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-76,114,-75.5</points>
<connection>
<GID>43</GID>
<name>IN_2</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112.5,-75.5,114,-75.5</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>114 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>112.5,-77.5,114,-77.5</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>114 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>114,-77.5,114,-77</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>-77.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133.5,-73.5,133.5,-72.5</points>
<connection>
<GID>45</GID>
<name>IN_7</name></connection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127.5,-72.5,133.5,-72.5</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<intersection>133.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,-74.5,133.5,-74.5</points>
<connection>
<GID>45</GID>
<name>IN_6</name></connection>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,-75.5,133.5,-75.5</points>
<connection>
<GID>45</GID>
<name>IN_5</name></connection>
<intersection>127.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>127.5,-76.5,127.5,-75.5</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>-75.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-77,133,-76.5</points>
<intersection>-77 2</intersection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-76.5,133.5,-76.5</points>
<connection>
<GID>45</GID>
<name>IN_4</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127.5,-77,133,-77</points>
<intersection>127.5 3</intersection>
<intersection>133 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>127.5,-78.5,127.5,-77</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>-77 2</intersection></vsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,-80.5,128,-77.5</points>
<intersection>-80.5 2</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128,-77.5,133.5,-77.5</points>
<connection>
<GID>45</GID>
<name>IN_3</name></connection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127.5,-80.5,128,-80.5</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>128 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,-82.5,129,-80</points>
<intersection>-82.5 2</intersection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129,-80,133.5,-80</points>
<intersection>129 0</intersection>
<intersection>133.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127.5,-82.5,129,-82.5</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<intersection>129 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>133.5,-80,133.5,-78.5</points>
<connection>
<GID>45</GID>
<name>IN_2</name></connection>
<intersection>-80 1</intersection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,-84.5,130.5,-79.5</points>
<intersection>-84.5 2</intersection>
<intersection>-79.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130.5,-79.5,133.5,-79.5</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127.5,-84.5,130.5,-84.5</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>130.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,-86.5,131.5,-80.5</points>
<intersection>-86.5 2</intersection>
<intersection>-80.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131.5,-80.5,133.5,-80.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>131.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127.5,-86.5,131.5,-86.5</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<intersection>131.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-101,115.5,-94</points>
<intersection>-101 7</intersection>
<intersection>-97 8</intersection>
<intersection>-95 19</intersection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>115.5,-94,136,-94</points>
<intersection>115.5 0</intersection>
<intersection>125 6</intersection>
<intersection>136 13</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>125,-101,125,-94</points>
<intersection>-101 10</intersection>
<intersection>-97 15</intersection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>115.5,-101,117,-101</points>
<connection>
<GID>69</GID>
<name>K</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>115.5,-97,117,-97</points>
<connection>
<GID>69</GID>
<name>J</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>125,-101,128,-101</points>
<connection>
<GID>70</GID>
<name>K</name></connection>
<intersection>125 6</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>136,-101,136,-94</points>
<intersection>-101 17</intersection>
<intersection>-97 18</intersection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>125,-97,128,-97</points>
<connection>
<GID>70</GID>
<name>J</name></connection>
<intersection>125 6</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>136,-101,138,-101</points>
<connection>
<GID>71</GID>
<name>K</name></connection>
<intersection>136 13</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>136,-97,138,-97</points>
<connection>
<GID>71</GID>
<name>J</name></connection>
<intersection>136 13</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>110,-95,115.5,-95</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,-101,124,-99</points>
<intersection>-101 2</intersection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124,-99,128,-99</points>
<connection>
<GID>70</GID>
<name>clock</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>123,-101,124,-101</points>
<connection>
<GID>69</GID>
<name>nQ</name></connection>
<intersection>124 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-101,135,-99</points>
<intersection>-101 2</intersection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-99,138,-99</points>
<connection>
<GID>71</GID>
<name>clock</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>134,-101,135,-101</points>
<connection>
<GID>70</GID>
<name>nQ</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>145,-107,145,-97</points>
<intersection>-107 5</intersection>
<intersection>-97 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>144,-97,145,-97</points>
<connection>
<GID>71</GID>
<name>Q</name></connection>
<intersection>145 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>145,-107,150.5,-107</points>
<intersection>145 3</intersection>
<intersection>150.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>150.5,-107,150.5,-100.5</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>-107 5</intersection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-104.5,123.5,-97</points>
<intersection>-104.5 2</intersection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-97,123.5,-97</points>
<connection>
<GID>69</GID>
<name>Q</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>123.5,-104.5,147,-104.5</points>
<intersection>123.5 0</intersection>
<intersection>147 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>147,-104.5,147,-98.5</points>
<intersection>-104.5 2</intersection>
<intersection>-98.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>147,-98.5,150.5,-98.5</points>
<connection>
<GID>75</GID>
<name>IN_2</name></connection>
<intersection>147 4</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134.5,-106,134.5,-97</points>
<intersection>-106 3</intersection>
<intersection>-97 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>134.5,-106,148,-106</points>
<intersection>134.5 0</intersection>
<intersection>148 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>148,-106,148,-99.5</points>
<intersection>-106 3</intersection>
<intersection>-99.5 7</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>134,-97,134.5,-97</points>
<connection>
<GID>70</GID>
<name>Q</name></connection>
<intersection>134.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>148,-99.5,150.5,-99.5</points>
<connection>
<GID>75</GID>
<name>IN_1</name></connection>
<intersection>148 4</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>114.5,-99,117,-99</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>117 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>117,-99,117,-99</points>
<connection>
<GID>69</GID>
<name>clock</name></connection>
<intersection>-99 1</intersection></vsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>99.5,-99,100.5,-99</points>
<connection>
<GID>83</GID>
<name>CLK</name></connection>
<connection>
<GID>81</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-95,101.5,-95</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<connection>
<GID>85</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>115,-120,117.5,-120</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>117.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>117.5,-120,117.5,-120</points>
<connection>
<GID>91</GID>
<name>clock</name></connection>
<intersection>-120 1</intersection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>102,-120,103,-120</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<connection>
<GID>97</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124.5,-129,157,-129</points>
<connection>
<GID>103</GID>
<name>IN_2</name></connection>
<intersection>124.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>124.5,-129,124.5,-118</points>
<intersection>-129 1</intersection>
<intersection>-120 7</intersection>
<intersection>-118 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>123.5,-118,124.5,-118</points>
<connection>
<GID>91</GID>
<name>Q</name></connection>
<intersection>124.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>124.5,-120,128.5,-120</points>
<connection>
<GID>92</GID>
<name>clock</name></connection>
<intersection>124.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-132,135.5,-118</points>
<intersection>-132 1</intersection>
<intersection>-118 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-132,156,-132</points>
<intersection>135.5 0</intersection>
<intersection>136.5 4</intersection>
<intersection>156 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>134.5,-118,135.5,-118</points>
<connection>
<GID>92</GID>
<name>Q</name></connection>
<intersection>135.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>156,-132,156,-122</points>
<intersection>-132 1</intersection>
<intersection>-130 7</intersection>
<intersection>-122 6</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>136.5,-132,136.5,-120</points>
<intersection>-132 1</intersection>
<intersection>-120 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>136.5,-120,138.5,-120</points>
<connection>
<GID>93</GID>
<name>clock</name></connection>
<intersection>136.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>154,-122,156,-122</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>156 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>156,-130,157,-130</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>156 3</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,-131,148.5,-118</points>
<intersection>-131 2</intersection>
<intersection>-122 3</intersection>
<intersection>-118 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144.5,-118,148.5,-118</points>
<connection>
<GID>93</GID>
<name>Q</name></connection>
<intersection>148.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148.5,-131,157,-131</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>148.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>148.5,-122,152,-122</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>148.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153,-129.5,153,-128</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<intersection>-129.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>120.5,-129.5,120.5,-124</points>
<connection>
<GID>91</GID>
<name>clear</name></connection>
<intersection>-129.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>120.5,-129.5,153,-129.5</points>
<intersection>120.5 1</intersection>
<intersection>131.5 3</intersection>
<intersection>141.5 4</intersection>
<intersection>153 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>131.5,-129.5,131.5,-124</points>
<connection>
<GID>92</GID>
<name>clear</name></connection>
<intersection>-129.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>141.5,-129.5,141.5,-124</points>
<connection>
<GID>93</GID>
<name>clear</name></connection>
<intersection>-129.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-118,115,-116.5</points>
<intersection>-118 1</intersection>
<intersection>-116.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-118,117.5,-118</points>
<connection>
<GID>91</GID>
<name>J</name></connection>
<intersection>115 0</intersection>
<intersection>116 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>112.5,-116.5,115,-116.5</points>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>116,-122,116,-118</points>
<intersection>-122 4</intersection>
<intersection>-118 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>116,-122,117.5,-122</points>
<connection>
<GID>91</GID>
<name>K</name></connection>
<intersection>116 3</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,-122,127.5,-116</points>
<intersection>-122 4</intersection>
<intersection>-118 2</intersection>
<intersection>-116 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,-116,127.5,-116</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127.5,-118,128.5,-118</points>
<connection>
<GID>92</GID>
<name>J</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>127.5,-122,128.5,-122</points>
<connection>
<GID>92</GID>
<name>K</name></connection>
<intersection>127.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-122,138,-116</points>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection>
<intersection>-122 3</intersection>
<intersection>-118 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-118,138.5,-118</points>
<connection>
<GID>93</GID>
<name>J</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>138,-122,138.5,-122</points>
<connection>
<GID>93</GID>
<name>K</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>114.5,-149.5,117,-149.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>117 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>117,-149.5,117,-149.5</points>
<connection>
<GID>108</GID>
<name>clock</name></connection>
<intersection>-149.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>101.5,-149.5,102.5,-149.5</points>
<connection>
<GID>113</GID>
<name>CLK</name></connection>
<connection>
<GID>112</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152.5,-159,152.5,-157.5</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<intersection>-159 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>120,-159,120,-153.5</points>
<connection>
<GID>108</GID>
<name>clear</name></connection>
<intersection>-159 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>120,-159,152.5,-159</points>
<intersection>120 1</intersection>
<intersection>131 3</intersection>
<intersection>141 4</intersection>
<intersection>152.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>131,-159,131,-153.5</points>
<connection>
<GID>109</GID>
<name>clear</name></connection>
<intersection>-159 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>141,-159,141,-153.5</points>
<connection>
<GID>110</GID>
<name>clear</name></connection>
<intersection>-159 2</intersection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-151.5,115,-143</points>
<intersection>-151.5 2</intersection>
<intersection>-147.5 6</intersection>
<intersection>-143 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-143,136.5,-143</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection>
<intersection>126 4</intersection>
<intersection>136.5 11</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-151.5,117,-151.5</points>
<connection>
<GID>108</GID>
<name>K</name></connection>
<intersection>115 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>126,-151.5,126,-143</points>
<intersection>-151.5 9</intersection>
<intersection>-147.5 13</intersection>
<intersection>-143 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>115,-147.5,117,-147.5</points>
<connection>
<GID>108</GID>
<name>J</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>126,-151.5,128,-151.5</points>
<connection>
<GID>109</GID>
<name>K</name></connection>
<intersection>126 4</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>136.5,-151.5,136.5,-143</points>
<intersection>-151.5 15</intersection>
<intersection>-147.5 16</intersection>
<intersection>-143 1</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>126,-147.5,128,-147.5</points>
<connection>
<GID>109</GID>
<name>J</name></connection>
<intersection>126 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>136.5,-151.5,138,-151.5</points>
<connection>
<GID>110</GID>
<name>K</name></connection>
<intersection>136.5 11</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>136.5,-147.5,138,-147.5</points>
<connection>
<GID>110</GID>
<name>J</name></connection>
<intersection>136.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-143.5,99.5,-143.5</points>
<connection>
<GID>116</GID>
<name>OUT_0</name></connection>
<intersection>-143.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,-143.5,99.5,-143.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-149.5,124.5,-138.5</points>
<intersection>-149.5 1</intersection>
<intersection>-147.5 2</intersection>
<intersection>-138.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124.5,-149.5,128,-149.5</points>
<connection>
<GID>109</GID>
<name>clock</name></connection>
<intersection>124.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>123,-147.5,124.5,-147.5</points>
<connection>
<GID>108</GID>
<name>Q</name></connection>
<intersection>124.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>124.5,-138.5,127.5,-138.5</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>124.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-168,135,-144.5</points>
<intersection>-168 6</intersection>
<intersection>-149.5 5</intersection>
<intersection>-147.5 2</intersection>
<intersection>-144.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-144.5,153.5,-144.5</points>
<intersection>135 0</intersection>
<intersection>153.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>134,-147.5,135,-147.5</points>
<connection>
<GID>109</GID>
<name>Q</name></connection>
<intersection>135 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>153.5,-151.5,153.5,-144.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>-144.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>135,-149.5,138,-149.5</points>
<connection>
<GID>110</GID>
<name>clock</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>135,-168,137,-168</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145,-164.5,145,-147.5</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>-151.5 3</intersection>
<intersection>-147.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144,-147.5,145,-147.5</points>
<connection>
<GID>110</GID>
<name>Q</name></connection>
<intersection>145 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>145,-151.5,151.5,-151.5</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>145 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-160,160,-138.5</points>
<intersection>-160 1</intersection>
<intersection>-138.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160,-160,161.5,-160</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139,-138.5,160,-138.5</points>
<connection>
<GID>128</GID>
<name>N_in0</name></connection>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>160 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-168,151,-159.5</points>
<intersection>-168 2</intersection>
<intersection>-159.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-159.5,157,-159.5</points>
<intersection>151 0</intersection>
<intersection>157 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148.5,-168,151,-168</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<connection>
<GID>130</GID>
<name>N_in0</name></connection>
<intersection>151 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>157,-159.5,157,-159</points>
<intersection>-159.5 1</intersection>
<intersection>-159 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>157,-159,161.5,-159</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<intersection>157 3</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-164.5,156,-158</points>
<intersection>-164.5 2</intersection>
<intersection>-158 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156,-158,161.5,-158</points>
<connection>
<GID>115</GID>
<name>IN_2</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156,-164.5,156.5,-164.5</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<connection>
<GID>131</GID>
<name>N_in0</name></connection>
<intersection>156 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>114,-194.5,137.5,-194.5</points>
<intersection>114 6</intersection>
<intersection>124.5 5</intersection>
<intersection>137.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>137.5,-194.5,137.5,-189</points>
<intersection>-194.5 1</intersection>
<intersection>-189 17</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>124.5,-194.5,124.5,-188.5</points>
<intersection>-194.5 1</intersection>
<intersection>-188.5 18</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>114,-194.5,114,-188.5</points>
<intersection>-194.5 1</intersection>
<intersection>-188.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>113,-188.5,115.5,-188.5</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<connection>
<GID>135</GID>
<name>clock</name></connection>
<intersection>114 6</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>137.5,-189,143,-189</points>
<connection>
<GID>137</GID>
<name>clock</name></connection>
<intersection>137.5 4</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>124.5,-188.5,127.5,-188.5</points>
<connection>
<GID>136</GID>
<name>clock</name></connection>
<intersection>124.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-188.5,96.5,-188.5</points>
<connection>
<GID>145</GID>
<name>CLK</name></connection>
<connection>
<GID>141</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133.5,-186.5,133.5,-182.5</points>
<connection>
<GID>136</GID>
<name>Q</name></connection>
<intersection>-186.5 2</intersection>
<intersection>-182.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133.5,-182.5,134,-182.5</points>
<connection>
<GID>147</GID>
<name>IN_1</name></connection>
<intersection>133.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>133.5,-186.5,135,-186.5</points>
<intersection>133.5 0</intersection>
<intersection>135 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>135,-186.5,135,-185.5</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>-186.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-191,141,-181.5</points>
<intersection>-191 4</intersection>
<intersection>-187 2</intersection>
<intersection>-181.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140,-181.5,141,-181.5</points>
<connection>
<GID>147</GID>
<name>OUT</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>141,-187,143,-187</points>
<connection>
<GID>137</GID>
<name>J</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>141,-191,143,-191</points>
<connection>
<GID>137</GID>
<name>K</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-186.5,123,-180.5</points>
<intersection>-186.5 2</intersection>
<intersection>-183.5 6</intersection>
<intersection>-180.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-180.5,134,-180.5</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121.5,-186.5,127.5,-186.5</points>
<connection>
<GID>135</GID>
<name>Q</name></connection>
<connection>
<GID>136</GID>
<name>J</name></connection>
<intersection>123 0</intersection>
<intersection>125.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>125.5,-190.5,125.5,-186.5</points>
<intersection>-190.5 5</intersection>
<intersection>-186.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>125.5,-190.5,127.5,-190.5</points>
<connection>
<GID>136</GID>
<name>K</name></connection>
<intersection>125.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>123,-183.5,123.5,-183.5</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-190.5,113.5,-185</points>
<intersection>-190.5 1</intersection>
<intersection>-186.5 2</intersection>
<intersection>-185 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-190.5,115.5,-190.5</points>
<connection>
<GID>135</GID>
<name>K</name></connection>
<intersection>113.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-186.5,115.5,-186.5</points>
<connection>
<GID>135</GID>
<name>J</name></connection>
<intersection>113.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>112,-185,113.5,-185</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,-184,92,-184</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<connection>
<GID>149</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149,-187,149,-182.5</points>
<connection>
<GID>137</GID>
<name>Q</name></connection>
<intersection>-182.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149,-182.5,149.5,-182.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>149 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,-189,157.5,-189</points>
<connection>
<GID>158</GID>
<name>IN_2</name></connection>
<intersection>-189 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-189,157.5,-189</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,-191.5,157,-190</points>
<intersection>-191.5 2</intersection>
<intersection>-190 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157,-190,157.5,-190</points>
<connection>
<GID>158</GID>
<name>IN_1</name></connection>
<intersection>157 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-191.5,157,-191.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>157 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,-194.5,157.5,-191</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>-194.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-194.5,157.5,-194.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,30.9538,439.646,-233.338</PageViewport></page 1>
<page 2>
<PageViewport>0,30.9538,439.646,-233.338</PageViewport></page 2>
<page 3>
<PageViewport>0,30.9538,439.646,-233.338</PageViewport></page 3>
<page 4>
<PageViewport>0,30.9538,439.646,-233.338</PageViewport></page 4>
<page 5>
<PageViewport>0,30.9538,439.646,-233.338</PageViewport></page 5>
<page 6>
<PageViewport>0,30.9538,439.646,-233.338</PageViewport></page 6>
<page 7>
<PageViewport>0,30.9538,439.646,-233.338</PageViewport></page 7>
<page 8>
<PageViewport>0,30.9538,439.646,-233.338</PageViewport></page 8>
<page 9>
<PageViewport>0,30.9538,439.646,-233.338</PageViewport></page 9></circuit>